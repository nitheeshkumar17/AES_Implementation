module sub_bytes (
	input [7:0] text,
	output reg [7:0] sub_text);

always @(*) begin
case (text)
8'h01 : sub_text <= 8'h7C;
8'h02 : sub_text <= 8'h77;
8'h03 : sub_text <= 8'h7B;
8'h04 : sub_text <= 8'hF2;
8'h05 : sub_text <= 8'h6B;
8'h06 : sub_text <= 8'h6F;
8'h07 : sub_text <= 8'hC5;
8'h08 : sub_text <= 8'h30;
8'h09 : sub_text <= 8'h01;
8'h0A : sub_text <= 8'h67;
8'h0B : sub_text <= 8'h2B;
8'h0C : sub_text <= 8'hFE;
8'h0D : sub_text <= 8'hD7;
8'h0E : sub_text <= 8'hAB;
8'h0F : sub_text <= 8'h76;
8'h10 : sub_text <= 8'hCA;
8'h11 : sub_text <= 8'h82;
8'h12 : sub_text <= 8'hC9;
8'h13 : sub_text <= 8'h7D;
8'h14 : sub_text <= 8'hFA;
8'h15 : sub_text <= 8'h59;
8'h16 : sub_text <= 8'h47;
8'h17 : sub_text <= 8'hF0;
8'h18 : sub_text <= 8'hAD;
8'h19 : sub_text <= 8'hD4;
8'h1A : sub_text <= 8'hA2;
8'h1B : sub_text <= 8'hAF;
8'h1C : sub_text <= 8'h9C;
8'h1D : sub_text <= 8'hA4;
8'h1E : sub_text <= 8'h72;
8'h1F : sub_text <= 8'hC0;
8'h20 : sub_text <= 8'hB7;
8'h21 : sub_text <= 8'hFD;
8'h22 : sub_text <= 8'h93;
8'h23 : sub_text <= 8'h26;
8'h24 : sub_text <= 8'h36;
8'h25 : sub_text <= 8'h3F;
8'h26 : sub_text <= 8'hF7;
8'h27 : sub_text <= 8'hCC;
8'h28 : sub_text <= 8'h34;
8'h29 : sub_text <= 8'hA5;
8'h2A : sub_text <= 8'hE5;
8'h2B : sub_text <= 8'hF1;
8'h2C : sub_text <= 8'h71;
8'h2D : sub_text <= 8'hD8;
8'h2E : sub_text <= 8'h31;
8'h2F : sub_text <= 8'h15;
8'h30 : sub_text <= 8'h04;
8'h31 : sub_text <= 8'hC7;
8'h32 : sub_text <= 8'h23;
8'h33 : sub_text <= 8'hC3;
8'h34 : sub_text <= 8'h18;
8'h35 : sub_text <= 8'h96;
8'h36 : sub_text <= 8'h05;
8'h37 : sub_text <= 8'h9A;
8'h38 : sub_text <= 8'h07;
8'h39 : sub_text <= 8'h12;
8'h3A : sub_text <= 8'h80;
8'h3B : sub_text <= 8'hE2;
8'h3C : sub_text <= 8'hEB;
8'h3D : sub_text <= 8'h27;
8'h3E : sub_text <= 8'hB2;
8'h3F : sub_text <= 8'h75;
8'h40 : sub_text <= 8'h09;
8'h41 : sub_text <= 8'h83;
8'h42 : sub_text <= 8'h2C;
8'h43 : sub_text <= 8'h1A;
8'h44 : sub_text <= 8'h1B;
8'h45 : sub_text <= 8'h6E;
8'h46 : sub_text <= 8'h5A;
8'h47 : sub_text <= 8'hA0;
8'h48 : sub_text <= 8'h52;
8'h49 : sub_text <= 8'h3B;
8'h4A : sub_text <= 8'hD6;
8'h4B : sub_text <= 8'hB3;
8'h4C : sub_text <= 8'h29;
8'h4D : sub_text <= 8'hE3;
8'h4E : sub_text <= 8'h2F;
8'h4F : sub_text <= 8'h84;
8'h50 : sub_text <= 8'h53;
8'h51 : sub_text <= 8'hD1;
8'h52 : sub_text <= 8'h00;
8'h53 : sub_text <= 8'hED;
8'h54 : sub_text <= 8'h20;
8'h55 : sub_text <= 8'hFC;
8'h56 : sub_text <= 8'hB1;
8'h57 : sub_text <= 8'h5B;
8'h58 : sub_text <= 8'h6A;
8'h59 : sub_text <= 8'hCB;
8'h5A : sub_text <= 8'hBE;
8'h5B : sub_text <= 8'h39;
8'h5C : sub_text <= 8'h4A;
8'h5D : sub_text <= 8'h4C;
8'h5E : sub_text <= 8'h58;
8'h5F : sub_text <= 8'hCF;
8'h60 : sub_text <= 8'hD0;
8'h61 : sub_text <= 8'hEF;
8'h62 : sub_text <= 8'hAA;
8'h63 : sub_text <= 8'hFB;
8'h64 : sub_text <= 8'h43;
8'h65 : sub_text <= 8'h4D;
8'h66 : sub_text <= 8'h33;
8'h67 : sub_text <= 8'h85;
8'h68 : sub_text <= 8'h45;
8'h69 : sub_text <= 8'hF9;
8'h6A : sub_text <= 8'h02;
8'h6B : sub_text <= 8'h7F;
8'h6C : sub_text <= 8'h50;
8'h6D : sub_text <= 8'h3C;
8'h6E : sub_text <= 8'h9F;
8'h6F : sub_text <= 8'hA8;
8'h70 : sub_text <= 8'h51;
8'h71 : sub_text <= 8'hA3;
8'h72 : sub_text <= 8'h40;
8'h73 : sub_text <= 8'h8F;
8'h74 : sub_text <= 8'h92;
8'h75 : sub_text <= 8'h9D;
8'h76 : sub_text <= 8'h38;
8'h77 : sub_text <= 8'hF5;
8'h78 : sub_text <= 8'hBC;
8'h79 : sub_text <= 8'hB6;
8'h7A : sub_text <= 8'hDA;
8'h7B : sub_text <= 8'h21;
8'h7C : sub_text <= 8'h10;
8'h7D : sub_text <= 8'hFF;
8'h7E : sub_text <= 8'hF3;
8'h7F : sub_text <= 8'hD2;
8'h80 : sub_text <= 8'hCD;
8'h81 : sub_text <= 8'h0C;
8'h82 : sub_text <= 8'h13;
8'h83 : sub_text <= 8'hEC;
8'h84 : sub_text <= 8'h5F;
8'h85 : sub_text <= 8'h97;
8'h86 : sub_text <= 8'h44;
8'h87 : sub_text <= 8'h17;
8'h88 : sub_text <= 8'hC4;
8'h89 : sub_text <= 8'hA7;
8'h8A : sub_text <= 8'h7E;
8'h8B : sub_text <= 8'h3D;
8'h8C : sub_text <= 8'h64;
8'h8D : sub_text <= 8'h5D;
8'h8E : sub_text <= 8'h19;
8'h8F : sub_text <= 8'h73;
8'h90 : sub_text <= 8'h60;
8'h91 : sub_text <= 8'h81;
8'h92 : sub_text <= 8'h4F;
8'h93 : sub_text <= 8'hDC;
8'h94 : sub_text <= 8'h22;
8'h95 : sub_text <= 8'h2A;
8'h96 : sub_text <= 8'h90;
8'h97 : sub_text <= 8'h88;
8'h98 : sub_text <= 8'h46;
8'h99 : sub_text <= 8'hEE;
8'h9A : sub_text <= 8'hB8;
8'h9B : sub_text <= 8'h14;
8'h9C : sub_text <= 8'hDE;
8'h9D : sub_text <= 8'h5E;
8'h9E : sub_text <= 8'h0B;
8'h9F : sub_text <= 8'hDB;
8'hA0 : sub_text <= 8'hE0;
8'hA1 : sub_text <= 8'h32;
8'hA2 : sub_text <= 8'h3A;
8'hA3 : sub_text <= 8'h0A;
8'hA4 : sub_text <= 8'h49;
8'hA5 : sub_text <= 8'h06;
8'hA6 : sub_text <= 8'h24;
8'hA7 : sub_text <= 8'h5C;
8'hA8 : sub_text <= 8'hC2;
8'hA9 : sub_text <= 8'hD3;
8'hAA : sub_text <= 8'hAC;
8'hAB : sub_text <= 8'h62;
8'hAC : sub_text <= 8'h91;
8'hAD : sub_text <= 8'h95;
8'hAE : sub_text <= 8'hE4;
8'hAF : sub_text <= 8'h79;
8'hB0 : sub_text <= 8'hE7;
8'hB1 : sub_text <= 8'hC8;
8'hB2 : sub_text <= 8'h37;
8'hB3 : sub_text <= 8'h6D;
8'hB4 : sub_text <= 8'h8D;
8'hB5 : sub_text <= 8'hD5;
8'hB6 : sub_text <= 8'h4E;
8'hB7 : sub_text <= 8'hA9;
8'hB8 : sub_text <= 8'h6C;
8'hB9 : sub_text <= 8'h56;
8'hBA : sub_text <= 8'hF4;
8'hBB : sub_text <= 8'hEA;
8'hBC : sub_text <= 8'h65;
8'hBD : sub_text <= 8'h7A;
8'hBE : sub_text <= 8'hAE;
8'hBF : sub_text <= 8'h08;
8'hC0 : sub_text <= 8'hBA;
8'hC1 : sub_text <= 8'h78;
8'hC2 : sub_text <= 8'h25;
8'hC3 : sub_text <= 8'h2E;
8'hC4 : sub_text <= 8'h1C;
8'hC5 : sub_text <= 8'hA6;
8'hC6 : sub_text <= 8'hB4;
8'hC7 : sub_text <= 8'hC6;
8'hC8 : sub_text <= 8'hE8;
8'hC9 : sub_text <= 8'hDD;
8'hCA : sub_text <= 8'h74;
8'hCB : sub_text <= 8'h1F;
8'hCC : sub_text <= 8'h4B;
8'hCD : sub_text <= 8'hBD;
8'hCE : sub_text <= 8'h8B;
8'hCF : sub_text <= 8'h8A;
8'hD0 : sub_text <= 8'h70;
8'hD1 : sub_text <= 8'h3E;
8'hD2 : sub_text <= 8'hB5;
8'hD3 : sub_text <= 8'h66;
8'hD4 : sub_text <= 8'h48;
8'hD5 : sub_text <= 8'h03;
8'hD6 : sub_text <= 8'hF6;
8'hD7 : sub_text <= 8'h0E;
8'hD8 : sub_text <= 8'h61;
8'hD9 : sub_text <= 8'h35;
8'hDA : sub_text <= 8'h57;
8'hDB : sub_text <= 8'hB9;
8'hDC : sub_text <= 8'h86;
8'hDD : sub_text <= 8'hC1;
8'hDE : sub_text <= 8'h1D;
8'hDF : sub_text <= 8'h9E;
8'hE0 : sub_text <= 8'hE1;
8'hE1 : sub_text <= 8'hF8;
8'hE2 : sub_text <= 8'h98;
8'hE3 : sub_text <= 8'h11;
8'hE4 : sub_text <= 8'h69;
8'hE5 : sub_text <= 8'hD9;
8'hE6 : sub_text <= 8'h8E;
8'hE7 : sub_text <= 8'h94;
8'hE8 : sub_text <= 8'h9B;
8'hE9 : sub_text <= 8'h1E;
8'hEA : sub_text <= 8'h87;
8'hEB : sub_text <= 8'hE9;
8'hEC : sub_text <= 8'hCE;
8'hED : sub_text <= 8'h55;
8'hEE : sub_text <= 8'h28;
8'hEF : sub_text <= 8'hDF;
8'hF0 : sub_text <= 8'h8C;
8'hF1 : sub_text <= 8'hA1;
8'hF2 : sub_text <= 8'h89;
8'hF3 : sub_text <= 8'h0D;
8'hF4 : sub_text <= 8'hBF;
8'hF5 : sub_text <= 8'hE6;
8'hF6 : sub_text <= 8'h42;
8'hF7 : sub_text <= 8'h68;
8'hF8 : sub_text <= 8'h41;
8'hF9 : sub_text <= 8'h99;
8'hFA : sub_text <= 8'h2D;
8'hFB : sub_text <= 8'h0F;
8'hFC : sub_text <= 8'hB0;
8'hFD : sub_text <= 8'h54;
8'hFE : sub_text <= 8'hBB;
8'hFF : sub_text <= 8'h16;
default : sub_text <= 8'h00;
endcase
end 
endmodule
